/**
 *
 * Name:
 *   bp_fpga_host_io_in.sv
 *
 * Description:
 *   FPGA Host IO Input module with UART Rx from PC Host and io_cmd/resp to BP
 *
 * Inputs:
 *   io_resp_i - response to io_cmd_o messages
 *             - generate NBF packet to forward to bp_fpga_host_io_out
 *             - NBF packets generated include read reply, nbf fence done, nbf finish done
 *
 * Outputs:
 *   io_cmd_o - IO commands to BlackParrot generated from PC Host NBF packets
 *            - includes write and read memory, nbf fence, nbf finish
 *            - io_cmd_o may block if network is full
 *            - if backpressure builds and results in full NBF buffer and SIPO an RX
 *              error will be generated and forward to PC Host through bp_fpga_host_io_out
 *            - required throughput is determined by UART Baud Rate
 *            - with Baud Rate = 9600, 10 bits per byte (1 start, 8 data, 1 stop), and
 *              14 bytes per NBF command, this unit needs to process ~69 NBF commands
 *              per second. At Baud Rate = 115200, processing rate is ~823 NBF cmd/sec.
 *              At 10 MHz clock, that is ~144k cycles per cmd at 9600 Baud or ~12k cycles
 *              per cmd at 115200 Baud.
 *
 *   nbf_o - NBF packets to bp_fpga_host_io_out
 *         - generated by FSM processing io_resp_i, SIPO full enqueue error, and UART RX error
 *         - includes nbf finish, nbf fence done, UART RX error, memory read response
 *
 *
 * TODO:
 * NBF SIPO (bsg_serial_in_parallel_out_passthrough)
 * - convert UART RX bytes to NBF packet
 * - 1 byte input from UART RX to NBF packet (14 byte) output to NBF Buffer
 *
 * NBF Buffer (bsg_two_fifo or bsg_fifo_1r1w_small)
 * - buffer NBF packets from NBF SIPO
 *
 * Arbitration (bsg_arb_fixed)
 * - three inputs: io_resp_i FSM, SIPO enqueue error, UART RX error
 * - priority (high to low) = UART RX error, SIPO enqueue error, io_resp_i FSM
 * - outputs NBF packet on nbf_o port to bp_fpga_host_io_out
 *
 * FSM
 * - send io_cmd_o based on received NBF packets in NBF buffer
 * - sending should be non-blocking with processing io_resp_i so we don't stall the
 *   FSM and prevent it from consuming NBF buffer packets if io_cmd_o is available
 * - process io_resp_i and generate NBF packets for responses to PC Host - send to arbitration
 * - process NBF packets not requiring io_cmd to be sent.
 *   These include nbf fence and nbf finish
 *
 * io_cmd/resp credit flow control (bsg_flow_counter)
 * - credit flow control for cmd/resp network
 * - used by FSM to process nbf fence commands
 *
 */

module bp_fpga_host_io_in
  import bp_common_pkg::*;
  import bp_me_pkg::*;

  #(parameter bp_params_e bp_params_p = e_bp_default_cfg
    `declare_bp_proc_params(bp_params_p)

    , parameter nbf_addr_width_p = paddr_width_p
    , parameter nbf_data_width_p = dword_width_gp
    , localparam nbf_width_lp = `bp_fpga_host_nbf_width(nbf_addr_width_p, nbf_data_width_p)

    , parameter uart_clk_per_bit_p = 10416 // 100 MHz clock / 9600 Baud
    , parameter uart_data_bits_p = 8 // between 5 and 9 bits
    , parameter uart_parity_bit_p = 0 // 0 or 1
    , parameter uart_stop_bits_p = 1 // 1 or 2

    , parameter nbf_buffer_els_p = 4

    , localparam nbf_uart_packets_lp = (nbf_width_lp / uart_data_bits_p)

    `declare_bp_bedrock_mem_if_widths(paddr_width_p, cce_block_width_p, lce_id_width_p, lce_assoc_p, io)
    )
  (input                                     clk_i
   , input                                   reset_i

   // To BlackParrot
   , output logic [io_mem_msg_width_lp-1:0]  io_cmd_o
   , output logic                            io_cmd_v_o
   , input                                   io_cmd_yumi_i

   , input  [io_mem_msg_width_lp-1:0]        io_resp_i
   , input                                   io_resp_v_i
   , output logic                            io_resp_ready_and_o

   // UART to PC Host
   , input                                   rx_i

   // Signals to FPGA Host IO Out
   , output logic [nbf_width_lp-1:0]         nbf_o
   , output logic                            nbf_v_o
   , input                                   nbf_ready_and_i
   );

  `declare_bp_fpga_host_nbf_s(nbf_addr_width_p, nbf_data_width_p);

  logic rx_v_lo, rx_error_lo;
  logic [uart_data_bits_p-1:0] rx_data_lo;
  uart_rx
   #(.clk_per_bit_p(uart_clk_per_bit_p)
     ,.data_bits_p(uart_data_bits_p)
     ,.parity_bit_p(uart_parity_bit_p)
     ,.stop_bits_p(uart_stop_bits_p)
     )
    rx
    (.clk_i(clk_i)
     ,.reset_i(reset_i)
     ,.rx_i(rx_i)
     ,.rx_v_o(rx_v_lo)
     ,.rx_o(rx_data_lo)
     ,.rx_error_o(rx_error_lo)
     );

  logic nbf_sipo_ready_and_lo;
  logic nbf_sipo_v_lo, nbf_sipo_ready_and_li;
  bp_fpga_host_nbf_s nbf_lo;

  bsg_serial_in_parallel_out_passthrough
   #(.width_p(uart_data_bits_p)
     ,.els_p(nbf_uart_packets_lp)
     ,.hi_to_lo_p(0) // TODO: check this is correct order
     // byte order sent across UART RX should result in SIPO producing proper
     // NBF packet. UART RX will receive opcode byte, followed by LSB to MSB of
     // address then LSB to MSB of data
     )
    nbf_sipo
    (.clk_i(clk_i)
     ,.reset_i(reset_i)
     ,.v_i(rx_v_lo)
     ,.ready_and_o(nbf_sipo_ready_and_lo)
     ,.data_i(rx_data_lo)
     ,.data_o(nbf_lo)
     ,.v_o(nbf_sipo_v_lo)
     ,.ready_and_i(nbf_sipo_ready_and_li)
     );

  logic nbf_buffer_v_lo, nbf_buffer_yumi_li;
  bp_fpga_host_nbf_s nbf_buffer_lo;

  bsg_fifo_1r1w_small
   #(.width_p(nbf_width_lp)
     ,.els_p(nbf_buffer_els_p)
     ,.ready_THEN_valid_p(0)
     )
    nbf_fifo
    (.clk_i(clk_i)
     ,.reset_i(reset_i)
     ,.v_i(nbf_sipo_v_lo)
     ,.ready_o(nbf_sipo_ready_and_li)
     ,.data_i(nbf_lo)
     ,.v_o(nbf_buffer_v_lo)
     ,.data_o(nbf_buffer_lo)
     ,.yumi_i(nbf_buffer_yumi_li)
     );

  typedef enum logic [3:0]
  {

  } state_e;

  wire [2:0] arb_reqs_li = {rx_error_lo, nbf_sipo_error, io_nbf_v};
  logic [2:0] arb_grants_lo;
  bsg_arb_fixed
   #(.inputs_p(3)
     // order arb high to low
     ,.lo_to_hi_p(0)
     )
    nbf_out_arb
    (.ready_i(nbf_ready_and_i) // TODO: is this really a ready_then_v input?
     ,.reqs_i(arb_reqs_li)
     ,.grants_o(arb_grants_lo)
     );

  always_ff @(posedge clk_i) begin
  end

  always_comb begin
  end
 
endmodule
