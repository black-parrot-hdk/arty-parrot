/**
 *
 * Name:
 *   bp_fpga_host_io_in.sv
 *
 * Description:
 *   FPGA Host IO Input module with UART Rx from PC Host and io_cmd/resp to BP
 *
 * Inputs:
 *   io_resp_i - response to io_cmd_o messages
 *             - generate NBF packet to forward to bp_fpga_host_io_out
 *             - NBF packets generated include read reply, nbf fence done, nbf finish done
 *
 * Outputs:
 *   io_cmd_o - IO commands to BlackParrot generated from PC Host NBF packets
 *            - includes write and read memory, nbf fence, nbf finish
 *            - io_cmd_o may block if network is full
 *            - if backpressure builds and results in full NBF buffer and SIPO an RX
 *              error will be generated and forward to PC Host through bp_fpga_host_io_out
 *            - required throughput is determined by UART Baud Rate
 *            - with Baud Rate = 9600, 10 bits per byte (1 start, 8 data, 1 stop), and
 *              14 bytes per NBF command, this unit needs to process ~69 NBF commands
 *              per second. At Baud Rate = 115200, processing rate is ~823 NBF cmd/sec.
 *              At 10 MHz clock, that is ~144k cycles per cmd at 9600 Baud or ~12k cycles
 *              per cmd at 115200 Baud.
 *
 *   nbf_o - NBF packets to bp_fpga_host_io_out
 *         - generated by FSM processing io_resp_i, SIPO full enqueue error, and UART RX error
 *         - includes nbf finish, nbf fence done, UART RX error, memory read response
 *
 *
 * TODO:
 * Send error to PC Host on SIPO enqueue error or rx_error_o raised
 *
 */

`include "bp_common_defines.svh"
`include "bp_me_defines.svh"
`include "bp_fpga_host_defines.svh"

module bp_fpga_host_io_in
  import bp_common_pkg::*;
  import bp_me_pkg::*;
  import bp_fpga_host_pkg::*;

  #(parameter bp_params_e bp_params_p = e_bp_default_cfg
    `declare_bp_proc_params(bp_params_p)

    , parameter nbf_addr_width_p = paddr_width_p
    , parameter nbf_data_width_p = dword_width_gp
    , localparam nbf_width_lp = `bp_fpga_host_nbf_width(nbf_addr_width_p, nbf_data_width_p)

    , parameter uart_clk_per_bit_p = 10416 // 100 MHz clock / 9600 Baud
    , parameter uart_data_bits_p = 8 // between 5 and 9 bits
    , parameter uart_parity_bit_p = 0 // 0 or 1
    , parameter uart_stop_bits_p = 1 // 1 or 2

    , parameter nbf_buffer_els_p = 4

    , localparam nbf_uart_packets_lp = (nbf_width_lp / uart_data_bits_p)

    `declare_bp_bedrock_mem_if_widths(paddr_width_p, cce_block_width_p, lce_id_width_p, lce_assoc_p, io)
    )
  (input                                     clk_i
   , input                                   reset_i

   // To BlackParrot
   , output logic [io_mem_msg_width_lp-1:0]  io_cmd_o
   , output logic                            io_cmd_v_o
   , input                                   io_cmd_yumi_i

   , input  [io_mem_msg_width_lp-1:0]        io_resp_i
   , input                                   io_resp_v_i
   , output logic                            io_resp_ready_and_o

   // UART to PC Host
   , input                                   rx_i

   // Signals to FPGA Host IO Out
   , output logic [nbf_width_lp-1:0]         nbf_o
   , output logic                            nbf_v_o
   , input                                   nbf_ready_and_i

   // Error signal for debug
   // - implemented as a sticky bit
   , output logic                            error_o
   );

  `declare_bp_bedrock_mem_if(paddr_width_p, cce_block_width_p, lce_id_width_p, lce_assoc_p, io)
  `declare_bp_fpga_host_nbf_s(nbf_addr_width_p, nbf_data_width_p);

  bp_bedrock_io_mem_msg_s io_cmd, io_resp;
  assign io_cmd_o = io_cmd;
  bp_bedrock_io_mem_msg_payload_s io_cmd_payload;

  logic io_resp_v_lo, io_resp_yumi_li;
  // IO response buffer
  bsg_two_fifo
   #(.width_p($bits(bp_bedrock_io_mem_msg_s)))
    io_resp_fifo
     (.clk_i(clk_i)
      ,.reset_i(reset_i)
      // from input
      ,.v_i(io_resp_v_i)
      ,.ready_o(io_resp_ready_and_o)
      ,.data_i(io_resp_i)
      // to FSM
      ,.v_o(io_resp_v_lo)
      ,.yumi_i(io_resp_yumi_li)
      ,.data_o(io_resp)
      );


  bp_fpga_host_nbf_s nbf_lo;
  assign nbf_o = nbf_lo;

  logic rx_v_lo, rx_error_lo;
  logic [uart_data_bits_p-1:0] rx_data_lo;
  uart_rx
   #(.clk_per_bit_p(uart_clk_per_bit_p)
     ,.data_bits_p(uart_data_bits_p)
     ,.parity_bit_p(uart_parity_bit_p)
     ,.stop_bits_p(uart_stop_bits_p)
     )
    rx
    (.clk_i(clk_i)
     ,.reset_i(reset_i)
     // from PC / UART pin
     ,.rx_i(rx_i)
     // to nbf_sipo
     ,.rx_v_o(rx_v_lo)
     ,.rx_o(rx_data_lo)
     // error signal
     ,.rx_error_o(rx_error_lo)
     );

  logic nbf_sipo_ready_and_lo;
  logic nbf_sipo_v_lo, nbf_sipo_ready_and_li;
  bp_fpga_host_nbf_s nbf_sipo_lo;

  // Process bytes from UART RX
  // NBF packet arrives opcode, address (LSB to MSB), data (LSB to MSB)
  bsg_serial_in_parallel_out_passthrough
   #(.width_p(uart_data_bits_p)
     ,.els_p(nbf_uart_packets_lp)
     ,.hi_to_lo_p(0)
     )
    nbf_sipo
    (.clk_i(clk_i)
     ,.reset_i(reset_i)
     // from UART RX
     ,.v_i(rx_v_lo)
     ,.ready_and_o(nbf_sipo_ready_and_lo)
     ,.data_i(rx_data_lo)
     // to nbf_buffer
     ,.v_o(nbf_sipo_v_lo)
     ,.ready_and_i(nbf_sipo_ready_and_li)
     ,.data_o(nbf_sipo_lo)
     );

  logic nbf_buffer_v_lo, nbf_buffer_yumi_li;
  bp_fpga_host_nbf_s nbf_buffer_lo;

  bsg_fifo_1r1w_small
   #(.width_p(nbf_width_lp)
     ,.els_p(nbf_buffer_els_p)
     ,.ready_THEN_valid_p(0)
     )
    nbf_buffer
    (.clk_i(clk_i)
     ,.reset_i(reset_i)
     // from nbf_sipo
     ,.v_i(nbf_sipo_v_lo)
     ,.ready_o(nbf_sipo_ready_and_li)
     ,.data_i(nbf_sipo_lo)
     // to FSM
     ,.v_o(nbf_buffer_v_lo)
     ,.yumi_i(nbf_buffer_yumi_li)
     ,.data_o(nbf_buffer_lo)
     );

  wire is_fence_packet = (nbf_buffer_lo.opcode == e_fpga_host_nbf_fence);
  wire is_finish_packet = (nbf_buffer_lo.opcode == e_fpga_host_nbf_finish);

  typedef enum logic [1:0]
  {
    e_reset
    , e_send_nbf
  } io_in_state_e;

  io_in_state_e state_r, state_n;

  logic [`BSG_WIDTH(io_noc_max_credits_p)-1:0] credit_count_lo;
  bsg_flow_counter
   #(.els_p(io_noc_max_credits_p))
   nbf_counter
    (.clk_i(clk_i)
     ,.reset_i(reset_i)
     ,.v_i(io_cmd_yumi_i)
     ,.ready_i(1'b1)
     ,.yumi_i(io_resp_yumi_li)
     ,.count_o(credit_count_lo)
     );
  wire credits_full_lo = (credit_count_lo == io_noc_max_credits_p);
  wire credits_empty_lo = (credit_count_lo == '0);

  // sticky error bit
  // sources are UART RX and enqueue to SIPO when not ready
  logic error_r, error_n;
  assign error_n = ~reset_i & (rx_error_lo | (rx_v_lo & ~nbf_sipo_ready_and_lo));
  assign error_o = error_r;

  always_ff @(posedge clk_i) begin
    if (reset_i) begin
      error_r <= 1'b0;
      state_r <= e_reset;
    end else begin
      error_r <= error_r | error_n;
      state_r <= state_n;
    end
  end

  // nbf buffer sends packet to nbf_o port for finish and fence
  wire nbf_buffer_to_nbf_o = nbf_buffer_v_lo & (is_finish_packet | (credits_empty_lo & is_fence_packet));

  always_comb begin

    // outputs
    nbf_lo = '0;
    nbf_v_o = '0;
    io_cmd_v_o = '0;
    io_cmd = '0;

    // bufer dequeue signals
    io_resp_yumi_li = 1'b0;
    nbf_buffer_yumi_li = '0;

    // form io_cmd from current nbf_buffer output
    io_cmd.data = {'0, nbf_buffer_lo.data};
    io_cmd_payload = '0;
    // TODO: why does bp_top testbench pass this to bp_nonsynth_nbf_loader as LCE ID?
    io_cmd_payload.lce_id = lce_id_width_p'('b10);
    io_cmd.header.payload = io_cmd_payload;
    io_cmd.header.addr = nbf_buffer_lo.addr;
    unique case (nbf_bufer_lo.opcode)
      e_fpga_host_nbf_write_4: begin
        io_cmd.header.size = e_bedrock_msg_size_4;
        io_cmd.header.msg_type.mem = e_bedrock_mem_uc_wr;
        io_cmd.header.subop = e_bedrock_store;
      end
      e_fpga_host_nbf_write_8: begin
        io_cmd.header.size = e_bedrock_msg_size_8;
        io_cmd.header.msg_type.mem = e_bedrock_mem_uc_wr;
        io_cmd.header.subop = e_bedrock_store;
      end
      e_fpga_host_nbf_read_4: begin
        io_cmd.header.size = e_bedrock_msg_size_4;
        io_cmd.header.msg_type.mem = e_bedrock_mem_uc_rd;
      end
      e_fpga_host_nbf_read_8: begin
        io_cmd.header.size = e_bedrock_msg_size_8;
        io_cmd.header.msg_type.mem = e_bedrock_mem_uc_rd;
      end
      default: begin end
    endcase

    unique case (state_r)
      e_reset: begin
        state_n = reset_i ? e_reset : e_send_nbf;
      end
      e_send_nbf: begin
        // Current NBF command from PC Host is in nbf_buffer - two options:
        // 1. send command to BlackParrot over io_cmd_o
        // 2. send NBF response back to PC Host through bp_fpga_host_io_out

        // IO Resp for reads may also try to send NBF response to PC Host
        // through bp_fpga_host_io_out, but have lower priority than NBF buffer

        // Option 1 - send io_cmd_o
        // send IO command for current NBF command
        // requires available credits and that NBF cmd is not fence or finish
        io_cmd_v_o = nbf_buffer_v_lo & ~credits_full_lo
                     & ~is_fence_packet & ~is_finish_packet;

        // Option 2 - send nbf_o back to PC Host
        // send NBF packet to bp_fpga_host_io_out for current NBF command
        // if required (fence or finish)
        nbf_v_o = nbf_buffer_to_nbf_o;
        if (is_fence_packet) begin
          nbf_lo.opcode = e_fpga_host_nbf_fence;
        end else if (is_finish_packet) begin
          nbf_lo.opcode = e_fpga_host_nbf_finish;
        end

        // consume current NBF command from buffer when it either sends
        // on IO network or handshakes with bp_fpga_host_io_out
        nbf_buffer_yumi_li = io_cmd_yumi_i | (nbf_v_o & nbf_ready_and_i);

        // Process IO responses
        if (io_resp_v_lo) begin
          unique case (io_resp.header.msg_type.mem)
            // uc_wr was NBF store to BP - sink response
            e_bedrock_mem_uc_wr: begin
              io_resp_yumi_li = 1'b1;
            end
            // uc_rd is response from NBF read from BP - send NBF packet
            // to bp_fpga_host_io_out
            e_bedrock_mem_uc_rd: begin
              // can only process if nbf_o not in use
              if (~nbf_buffer_to_nbf_o) begin
                nbf_v_o = 1'b1;
                io_resp_yumi_li = nbf_ready_and_i;
                unique case (io_resp.header.size)
                  e_bedrock_msg_size_4: nbf_lo.opcode = e_fpga_host_nbf_read_4;
                  e_bedrock_msg_size_8: nbf_lo.opcode = e_fpga_host_nbf_read_8;
                  default: nbf_lo.opcode = e_fpga_host_nbf_error;
                endcase
                nbf_lo.addr = io_resp.header.addr;
                nbf_lo.data = io_resp.data[0+:nbf_data_width_p];
              end
            end
            default: begin end
          endcase // io_resp msg_type
        end // io_resp_v_lo
      end // e_send_nbf
      default: begin end
    endcase // state_r
  end // always_comb
 
endmodule
