/*
 * bp_fpga_host_pkg.sv
 *
 * Contains the FPGA Host to PC Host NBF structures.
 *
 */

 package bp_fpga_host_pkg;

  `include "bp_fpga_host_pkgdef.svh"

 endpackage
