`ifndef uart_defs_vh
`define uart_defs_vh

`define SAFE_CLOG2(x) (((x)==1) ? 1 : $clog2((x)))

`endif